`timescale 1ns / 1ps
module FullAdder(
    input  wire a,
    input  wire b,
    input  wire cin,
    output wire sum,
    output wire cout
);
    assign sum  = a ^ b ^ cin; // bool expression for sum 
    assign cout = (a & b) | (b & cin) | (a & cin);
endmodule